--**********************************************
-- 	UNIVERSIDAD AUTONOMA DE SAN LUIS POTOSI  
-- 	School of Sciences                         
-- 	Author: Octavio Torres Delgado           
--**********************************************

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity learningRates is
	port( weight1 : in std_logic_vector(15 downto 0);
		  weight2 : in std_logic_vector(15 downto 0);
		  weight3 : in std_logic_vector(15 downto 0);  
  
		  nk1 : out std_logic_vector(4 downto 0);
		  nk2 : out std_logic_vector(4 downto 0);
		  nk3 : out std_logic_vector(4 downto 0));
end entity;

architecture learningRates_architecture of learningRates is

-- LUTs for the computing of log2(alpha_k,t) = log2(alphaw/wk,t)
-- alphaw = 0.001953125 = 2^⁻9
type memory is array (0 to 255) of std_logic_vector(4 downto 0);

CONSTANT log2_memory1 : memory :=
(
	0 => "11111", -- -1.0
    1 => "11111", -- -1.0
	2 => "11110", -- -2.0
    3 => "11101", -- -3.0
    4 => "11101", -- -3.0
    5 => "11101", -- -3.0
	6 => "11100", -- -4.0
	7 => "11100", -- -4.0
	8 => "11100", -- -4.0
	9 => "11100", -- -4.0
	10 => "11100", -- -4.0
	11 => "11100", -- -4.0
    12 => "11011", -- -5.0
    13 => "11011", -- -5.0
	14 => "11011", -- -5.0
	15 => "11011", -- -5.0
	16 => "11011", -- -5.0
	17 => "11011", -- -5.0
	18 => "11011", -- -5.0
	19 => "11011", -- -5.0
	20 => "11011", -- -5.0
	21 => "11011", -- -5.0
	22 => "11011", -- -5.0
	23 => "11010", -- -6.0
	24 => "11010", -- -6.0
	25 => "11010", -- -6.0
	26 => "11010", -- -6.0
	27 => "11010", -- -6.0
	28 => "11010", -- -6.0
	29 => "11010", -- -6.0
	30 => "11010", -- -6.0
	31 => "11010", -- -6.0
	32 => "11010", -- -6.0
	33 => "11010", -- -6.0
	34 => "11010", -- -6.0
	35 => "11010", -- -6.0
	36 => "11010", -- -6.0
	37 => "11010", -- -6.0
	38 => "11010", -- -6.0
	39 => "11010", -- -6.0
	40 => "11010", -- -6.0
	41 => "11010", -- -6.0
	42 => "11010", -- -6.0
	43 => "11010", -- -6.0
	44 => "11010", -- -6.0
	45 => "11010", -- -6.0
	46 => "11001", -- -7.0
	47 => "11001", -- -7.0
	48 => "11001", -- -7.0
	49 => "11001", -- -7.0
	50 => "11001", -- -7.0
	51 => "11001", -- -7.0
	52 => "11001", -- -7.0
	53 => "11001", -- -7.0
	54 => "11001", -- -7.0
	55 => "11001", -- -7.0
	56 => "11001", -- -7.0
	57 => "11001", -- -7.0
	58 => "11001", -- -7.0
	59 => "11001", -- -7.0
	60 => "11001", -- -7.0
	61 => "11001", -- -7.0
	62 => "11001", -- -7.0
	63 => "11001", -- -7.0
	64 => "11001", -- -7.0
	65 => "11001", -- -7.0
	66 => "11001", -- -7.0
	67 => "11001", -- -7.0
	68 => "11001", -- -7.0
	69 => "11001", -- -7.0
	70 => "11001", -- -7.0
	71 => "11001", -- -7.0
	72 => "11001", -- -7.0
	73 => "11001", -- -7.0
	74 => "11001", -- -7.0
	75 => "11001", -- -7.0
	76 => "11001", -- -7.0
	77 => "11001", -- -7.0
	78 => "11001", -- -7.0
	79 => "11001", -- -7.0
	80 => "11001", -- -7.0
	81 => "11001", -- -7.0
	82 => "11001", -- -7.0
	83 => "11001", -- -7.0
	84 => "11001", -- -7.0
	85 => "11001", -- -7.0
	86 => "11001", -- -7.0
	87 => "11001", -- -7.0
	88 => "11001", -- -7.0
	89 => "11001", -- -7.0
	90 => "11001", -- -7.0
	91 => "11000", -- -8.0
	92 => "11000", -- -8.0
	93 => "11000", -- -8.0
	94 => "11000", -- -8.0
	95 => "11000", -- -8.0
	96 => "11000", -- -8.0
	97 => "11000", -- -8.0
	98 => "11000", -- -8.0
	99 => "11000", -- -8.0
	100 => "11000", -- -8.0
	101 => "11000", -- -8.0
	102 => "11000", -- -8.0
	103 => "11000", -- -8.0
	104 => "11000", -- -8.0
	105 => "11000", -- -8.0
	106 => "11000", -- -8.0
	107 => "11000", -- -8.0
	108 => "11000", -- -8.0
	109 => "11000", -- -8.0
	110 => "11000", -- -8.0
	111 => "11000", -- -8.0
	112 => "11000", -- -8.0
	113 => "11000", -- -8.0
	114 => "11000", -- -8.0
	115 => "11000", -- -8.0
	116 => "11000", -- -8.0
	117 => "11000", -- -8.0
	118 => "11000", -- -8.0
	119 => "11000", -- -8.0
	120 => "11000", -- -8.0
	121 => "11000", -- -8.0
	122 => "11000", -- -8.0
	123 => "11000", -- -8.0
	124 => "11000", -- -8.0
	125 => "11000", -- -8.0
	126 => "11000", -- -8.0
	127 => "11000", -- -8.0
	128 => "11000", -- -8.0
	129 => "11000", -- -8.0
	130 => "11000", -- -8.0
	131 => "11000", -- -8.0
	132 => "11000", -- -8.0
	133 => "11000", -- -8.0
	134 => "11000", -- -8.0
	135 => "11000", -- -8.0
	136 => "11000", -- -8.0
	137 => "11000", -- -8.0
	138 => "11000", -- -8.0
	139 => "11000", -- -8.0
	140 => "11000", -- -8.0
	141 => "11000", -- -8.0
	142 => "11000", -- -8.0
	143 => "11000", -- -8.0
	144 => "11000", -- -8.0
	145 => "11000", -- -8.0
	146 => "11000", -- -8.0
	147 => "11000", -- -8.0
	148 => "11000", -- -8.0
	149 => "11000", -- -8.0
	150 => "11000", -- -8.0
	151 => "11000", -- -8.0
	152 => "11000", -- -8.0
	153 => "11000", -- -8.0
	154 => "11000", -- -8.0
	155 => "11000", -- -8.0
	156 => "11000", -- -8.0
	157 => "11000", -- -8.0
	158 => "11000", -- -8.0
	159 => "11000", -- -8.0
	160 => "11000", -- -8.0
	161 => "11000", -- -8.0
	162 => "11000", -- -8.0
	163 => "11000", -- -8.0
	164 => "11000", -- -8.0
	165 => "11000", -- -8.0
	166 => "11000", -- -8.0
	167 => "11000", -- -8.0
	168 => "11000", -- -8.0
	169 => "11000", -- -8.0
	170 => "11000", -- -8.0
	171 => "11000", -- -8.0
	172 => "11000", -- -8.0
	173 => "11000", -- -8.0
	174 => "11000", -- -8.0
	175 => "11000", -- -8.0
	176 => "11000", -- -8.0
	177 => "11000", -- -8.0
	178 => "11000", -- -8.0
	179 => "11000", -- -8.0
	180 => "11000", -- -8.0
	181 => "11000", -- -8.0
	others => "10111"); -- -9.0


CONSTANT log2_memory2 : memory :=
(
	0 => "11111", -- -1.0
    1 => "11111", -- -1.0
	2 => "11110", -- -2.0
    3 => "11101", -- -3.0
    4 => "11101", -- -3.0
    5 => "11101", -- -3.0
	6 => "11100", -- -4.0
	7 => "11100", -- -4.0
	8 => "11100", -- -4.0
	9 => "11100", -- -4.0
	10 => "11100", -- -4.0
	11 => "11100", -- -4.0
    12 => "11011", -- -5.0
    13 => "11011", -- -5.0
	14 => "11011", -- -5.0
	15 => "11011", -- -5.0
	16 => "11011", -- -5.0
	17 => "11011", -- -5.0
	18 => "11011", -- -5.0
	19 => "11011", -- -5.0
	20 => "11011", -- -5.0
	21 => "11011", -- -5.0
	22 => "11011", -- -5.0
	23 => "11010", -- -6.0
	24 => "11010", -- -6.0
	25 => "11010", -- -6.0
	26 => "11010", -- -6.0
	27 => "11010", -- -6.0
	28 => "11010", -- -6.0
	29 => "11010", -- -6.0
	30 => "11010", -- -6.0
	31 => "11010", -- -6.0
	32 => "11010", -- -6.0
	33 => "11010", -- -6.0
	34 => "11010", -- -6.0
	35 => "11010", -- -6.0
	36 => "11010", -- -6.0
	37 => "11010", -- -6.0
	38 => "11010", -- -6.0
	39 => "11010", -- -6.0
	40 => "11010", -- -6.0
	41 => "11010", -- -6.0
	42 => "11010", -- -6.0
	43 => "11010", -- -6.0
	44 => "11010", -- -6.0
	45 => "11010", -- -6.0
	46 => "11001", -- -7.0
	47 => "11001", -- -7.0
	48 => "11001", -- -7.0
	49 => "11001", -- -7.0
	50 => "11001", -- -7.0
	51 => "11001", -- -7.0
	52 => "11001", -- -7.0
	53 => "11001", -- -7.0
	54 => "11001", -- -7.0
	55 => "11001", -- -7.0
	56 => "11001", -- -7.0
	57 => "11001", -- -7.0
	58 => "11001", -- -7.0
	59 => "11001", -- -7.0
	60 => "11001", -- -7.0
	61 => "11001", -- -7.0
	62 => "11001", -- -7.0
	63 => "11001", -- -7.0
	64 => "11001", -- -7.0
	65 => "11001", -- -7.0
	66 => "11001", -- -7.0
	67 => "11001", -- -7.0
	68 => "11001", -- -7.0
	69 => "11001", -- -7.0
	70 => "11001", -- -7.0
	71 => "11001", -- -7.0
	72 => "11001", -- -7.0
	73 => "11001", -- -7.0
	74 => "11001", -- -7.0
	75 => "11001", -- -7.0
	76 => "11001", -- -7.0
	77 => "11001", -- -7.0
	78 => "11001", -- -7.0
	79 => "11001", -- -7.0
	80 => "11001", -- -7.0
	81 => "11001", -- -7.0
	82 => "11001", -- -7.0
	83 => "11001", -- -7.0
	84 => "11001", -- -7.0
	85 => "11001", -- -7.0
	86 => "11001", -- -7.0
	87 => "11001", -- -7.0
	88 => "11001", -- -7.0
	89 => "11001", -- -7.0
	90 => "11001", -- -7.0
	91 => "11000", -- -8.0
	92 => "11000", -- -8.0
	93 => "11000", -- -8.0
	94 => "11000", -- -8.0
	95 => "11000", -- -8.0
	96 => "11000", -- -8.0
	97 => "11000", -- -8.0
	98 => "11000", -- -8.0
	99 => "11000", -- -8.0
	100 => "11000", -- -8.0
	101 => "11000", -- -8.0
	102 => "11000", -- -8.0
	103 => "11000", -- -8.0
	104 => "11000", -- -8.0
	105 => "11000", -- -8.0
	106 => "11000", -- -8.0
	107 => "11000", -- -8.0
	108 => "11000", -- -8.0
	109 => "11000", -- -8.0
	110 => "11000", -- -8.0
	111 => "11000", -- -8.0
	112 => "11000", -- -8.0
	113 => "11000", -- -8.0
	114 => "11000", -- -8.0
	115 => "11000", -- -8.0
	116 => "11000", -- -8.0
	117 => "11000", -- -8.0
	118 => "11000", -- -8.0
	119 => "11000", -- -8.0
	120 => "11000", -- -8.0
	121 => "11000", -- -8.0
	122 => "11000", -- -8.0
	123 => "11000", -- -8.0
	124 => "11000", -- -8.0
	125 => "11000", -- -8.0
	126 => "11000", -- -8.0
	127 => "11000", -- -8.0
	128 => "11000", -- -8.0
	129 => "11000", -- -8.0
	130 => "11000", -- -8.0
	131 => "11000", -- -8.0
	132 => "11000", -- -8.0
	133 => "11000", -- -8.0
	134 => "11000", -- -8.0
	135 => "11000", -- -8.0
	136 => "11000", -- -8.0
	137 => "11000", -- -8.0
	138 => "11000", -- -8.0
	139 => "11000", -- -8.0
	140 => "11000", -- -8.0
	141 => "11000", -- -8.0
	142 => "11000", -- -8.0
	143 => "11000", -- -8.0
	144 => "11000", -- -8.0
	145 => "11000", -- -8.0
	146 => "11000", -- -8.0
	147 => "11000", -- -8.0
	148 => "11000", -- -8.0
	149 => "11000", -- -8.0
	150 => "11000", -- -8.0
	151 => "11000", -- -8.0
	152 => "11000", -- -8.0
	153 => "11000", -- -8.0
	154 => "11000", -- -8.0
	155 => "11000", -- -8.0
	156 => "11000", -- -8.0
	157 => "11000", -- -8.0
	158 => "11000", -- -8.0
	159 => "11000", -- -8.0
	160 => "11000", -- -8.0
	161 => "11000", -- -8.0
	162 => "11000", -- -8.0
	163 => "11000", -- -8.0
	164 => "11000", -- -8.0
	165 => "11000", -- -8.0
	166 => "11000", -- -8.0
	167 => "11000", -- -8.0
	168 => "11000", -- -8.0
	169 => "11000", -- -8.0
	170 => "11000", -- -8.0
	171 => "11000", -- -8.0
	172 => "11000", -- -8.0
	173 => "11000", -- -8.0
	174 => "11000", -- -8.0
	175 => "11000", -- -8.0
	176 => "11000", -- -8.0
	177 => "11000", -- -8.0
	178 => "11000", -- -8.0
	179 => "11000", -- -8.0
	180 => "11000", -- -8.0
	181 => "11000", -- -8.0
	others => "10111"); -- -9.0

  
CONSTANT log2_memory3 : memory :=
(
	0 => "11111", -- -1.0
    1 => "11111", -- -1.0
	2 => "11110", -- -2.0
    3 => "11101", -- -3.0
    4 => "11101", -- -3.0
    5 => "11101", -- -3.0
	6 => "11100", -- -4.0
	7 => "11100", -- -4.0
	8 => "11100", -- -4.0
	9 => "11100", -- -4.0
	10 => "11100", -- -4.0
	11 => "11100", -- -4.0
    12 => "11011", -- -5.0
    13 => "11011", -- -5.0
	14 => "11011", -- -5.0
	15 => "11011", -- -5.0
	16 => "11011", -- -5.0
	17 => "11011", -- -5.0
	18 => "11011", -- -5.0
	19 => "11011", -- -5.0
	20 => "11011", -- -5.0
	21 => "11011", -- -5.0
	22 => "11011", -- -5.0
	23 => "11010", -- -6.0
	24 => "11010", -- -6.0
	25 => "11010", -- -6.0
	26 => "11010", -- -6.0
	27 => "11010", -- -6.0
	28 => "11010", -- -6.0
	29 => "11010", -- -6.0
	30 => "11010", -- -6.0
	31 => "11010", -- -6.0
	32 => "11010", -- -6.0
	33 => "11010", -- -6.0
	34 => "11010", -- -6.0
	35 => "11010", -- -6.0
	36 => "11010", -- -6.0
	37 => "11010", -- -6.0
	38 => "11010", -- -6.0
	39 => "11010", -- -6.0
	40 => "11010", -- -6.0
	41 => "11010", -- -6.0
	42 => "11010", -- -6.0
	43 => "11010", -- -6.0
	44 => "11010", -- -6.0
	45 => "11010", -- -6.0
	46 => "11001", -- -7.0
	47 => "11001", -- -7.0
	48 => "11001", -- -7.0
	49 => "11001", -- -7.0
	50 => "11001", -- -7.0
	51 => "11001", -- -7.0
	52 => "11001", -- -7.0
	53 => "11001", -- -7.0
	54 => "11001", -- -7.0
	55 => "11001", -- -7.0
	56 => "11001", -- -7.0
	57 => "11001", -- -7.0
	58 => "11001", -- -7.0
	59 => "11001", -- -7.0
	60 => "11001", -- -7.0
	61 => "11001", -- -7.0
	62 => "11001", -- -7.0
	63 => "11001", -- -7.0
	64 => "11001", -- -7.0
	65 => "11001", -- -7.0
	66 => "11001", -- -7.0
	67 => "11001", -- -7.0
	68 => "11001", -- -7.0
	69 => "11001", -- -7.0
	70 => "11001", -- -7.0
	71 => "11001", -- -7.0
	72 => "11001", -- -7.0
	73 => "11001", -- -7.0
	74 => "11001", -- -7.0
	75 => "11001", -- -7.0
	76 => "11001", -- -7.0
	77 => "11001", -- -7.0
	78 => "11001", -- -7.0
	79 => "11001", -- -7.0
	80 => "11001", -- -7.0
	81 => "11001", -- -7.0
	82 => "11001", -- -7.0
	83 => "11001", -- -7.0
	84 => "11001", -- -7.0
	85 => "11001", -- -7.0
	86 => "11001", -- -7.0
	87 => "11001", -- -7.0
	88 => "11001", -- -7.0
	89 => "11001", -- -7.0
	90 => "11001", -- -7.0
	91 => "11000", -- -8.0
	92 => "11000", -- -8.0
	93 => "11000", -- -8.0
	94 => "11000", -- -8.0
	95 => "11000", -- -8.0
	96 => "11000", -- -8.0
	97 => "11000", -- -8.0
	98 => "11000", -- -8.0
	99 => "11000", -- -8.0
	100 => "11000", -- -8.0
	101 => "11000", -- -8.0
	102 => "11000", -- -8.0
	103 => "11000", -- -8.0
	104 => "11000", -- -8.0
	105 => "11000", -- -8.0
	106 => "11000", -- -8.0
	107 => "11000", -- -8.0
	108 => "11000", -- -8.0
	109 => "11000", -- -8.0
	110 => "11000", -- -8.0
	111 => "11000", -- -8.0
	112 => "11000", -- -8.0
	113 => "11000", -- -8.0
	114 => "11000", -- -8.0
	115 => "11000", -- -8.0
	116 => "11000", -- -8.0
	117 => "11000", -- -8.0
	118 => "11000", -- -8.0
	119 => "11000", -- -8.0
	120 => "11000", -- -8.0
	121 => "11000", -- -8.0
	122 => "11000", -- -8.0
	123 => "11000", -- -8.0
	124 => "11000", -- -8.0
	125 => "11000", -- -8.0
	126 => "11000", -- -8.0
	127 => "11000", -- -8.0
	128 => "11000", -- -8.0
	129 => "11000", -- -8.0
	130 => "11000", -- -8.0
	131 => "11000", -- -8.0
	132 => "11000", -- -8.0
	133 => "11000", -- -8.0
	134 => "11000", -- -8.0
	135 => "11000", -- -8.0
	136 => "11000", -- -8.0
	137 => "11000", -- -8.0
	138 => "11000", -- -8.0
	139 => "11000", -- -8.0
	140 => "11000", -- -8.0
	141 => "11000", -- -8.0
	142 => "11000", -- -8.0
	143 => "11000", -- -8.0
	144 => "11000", -- -8.0
	145 => "11000", -- -8.0
	146 => "11000", -- -8.0
	147 => "11000", -- -8.0
	148 => "11000", -- -8.0
	149 => "11000", -- -8.0
	150 => "11000", -- -8.0
	151 => "11000", -- -8.0
	152 => "11000", -- -8.0
	153 => "11000", -- -8.0
	154 => "11000", -- -8.0
	155 => "11000", -- -8.0
	156 => "11000", -- -8.0
	157 => "11000", -- -8.0
	158 => "11000", -- -8.0
	159 => "11000", -- -8.0
	160 => "11000", -- -8.0
	161 => "11000", -- -8.0
	162 => "11000", -- -8.0
	163 => "11000", -- -8.0
	164 => "11000", -- -8.0
	165 => "11000", -- -8.0
	166 => "11000", -- -8.0
	167 => "11000", -- -8.0
	168 => "11000", -- -8.0
	169 => "11000", -- -8.0
	170 => "11000", -- -8.0
	171 => "11000", -- -8.0
	172 => "11000", -- -8.0
	173 => "11000", -- -8.0
	174 => "11000", -- -8.0
	175 => "11000", -- -8.0
	176 => "11000", -- -8.0
	177 => "11000", -- -8.0
	178 => "11000", -- -8.0
	179 => "11000", -- -8.0
	180 => "11000", -- -8.0
	181 => "11000", -- -8.0
	others => "10111"); -- -9.0
  
begin
  
	-- Outputs  
  	nk1 <= log2_memory1(to_integer(unsigned(weight1(15 downto 8)))); 
  	nk2 <= log2_memory2(to_integer(unsigned(weight2(15 downto 8))));
  	nk3 <= log2_memory3(to_integer(unsigned(weight3(15 downto 8))));
    
end architecture;

